version https://git-lfs.github.com/spec/v1
oid sha256:e87a10b5672f54fb5085cbc1f305eb7057e741f8ddb32ff7c887c6ea2c7110ec
size 2152
